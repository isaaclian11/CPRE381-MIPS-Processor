-------------------------------------------------------------------------
-- Aidan Sherburne
-- Iowa State University
-------------------------------------------------------------------------
-- decoder_532_df.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: Dataflow 5:32 decoder for CPRE 381 Lab 3 P1e
-------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY decoder_532_df IS
  PORT (
    i_DecIn : IN std_logic_vector(4 DOWNTO 0); -- input binary encoded value
    o_DecOut : OUT std_logic_vector(31 DOWNTO 0)); -- output decoded bit

END decoder_532_df;
ARCHITECTURE dataflow OF decoder_532_df IS
BEGIN
  WITH i_DecIn SELECT o_DecOut <=

    "10000000000000000000000000000000" WHEN "11111",
    "01000000000000000000000000000000" WHEN "11110",
    "00100000000000000000000000000000" WHEN "11101",
    "00010000000000000000000000000000" WHEN "11100",
    "00001000000000000000000000000000" WHEN "11011",
    "00000100000000000000000000000000" WHEN "11010",
    "00000010000000000000000000000000" WHEN "11001",
    "00000001000000000000000000000000" WHEN "11000",
    "00000000100000000000000000000000" WHEN "10111",
    "00000000010000000000000000000000" WHEN "10110",
    "00000000001000000000000000000000" WHEN "10101",
    "00000000000100000000000000000000" WHEN "10100",
    "00000000000010000000000000000000" WHEN "10011",
    "00000000000001000000000000000000" WHEN "10010",
    "00000000000000100000000000000000" WHEN "10001",
    "00000000000000010000000000000000" WHEN "10000",
    "00000000000000001000000000000000" WHEN "01111",
    "00000000000000000100000000000000" WHEN "01110",
    "00000000000000000010000000000000" WHEN "01101",
    "00000000000000000001000000000000" WHEN "01100",
    "00000000000000000000100000000000" WHEN "01011",
    "00000000000000000000010000000000" WHEN "01010",
    "00000000000000000000001000000000" WHEN "01001",
    "00000000000000000000000100000000" WHEN "01000",
    "00000000000000000000000010000000" WHEN "00111",
    "00000000000000000000000001000000" WHEN "00110",
    "00000000000000000000000000100000" WHEN "00101",
    "00000000000000000000000000010000" WHEN "00100",
    "00000000000000000000000000001000" WHEN "00011",
    "00000000000000000000000000000100" WHEN "00010",
    "00000000000000000000000000000010" WHEN "00001",
    "00000000000000000000000000000001" WHEN "00000",
    "00000000000000000000000000000000" WHEN OTHERS;

END dataflow;